`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/29/2023 03:51:41 PM
// Design Name: 
// Module Name: game
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module game(
    input wire [1:0] mode,
    input wire CLK, // 100 Mhz clock
    input wire [7:0] keycode, // left and up buttons
    input wire [1:0] BTN_LU,
    input wire [1:0] BTN_DR,
    input wire switch,
    output wire VGA_HS, // horizontal sync
    output wire VGA_VS, // vertical sync
    output reg [3:0] VGA_R, // red channels
    output reg [3:0] VGA_G, // green channels
    output reg [3:0] VGA_B, // blue channels
    output wire [2:0] endgame, // game end flag
    output wire [8:0] lives1,lives2
    );
    
    wire lives1A,lives2A,lives10,lives20;
    
    localparam RW = 10; // rocket width
    localparam RH = 30; // rocket height
    localparam RY = 440 - RH; // initial paddle y
    localparam RX1 = 640-RW; // initial paddle x
    localparam RX = 0 + RW; // initial paddle x
    localparam RX3 = 320 - RW; // initial paddle x

    localparam IX = 300; // intial ball x
    localparam IY = 470 -RH - RH - 30; //initial ball y
    localparam IX2= 340;
    localparam B_SIZE = 10; // ball size
    localparam wall_l = 310;
    localparam wall_r = 330;
    localparam height = 477;
    
    reg [15:0] cnt = 0; // pixel clock counter
    reg pix_stb = 0; // pixel clock
    wire score;
    wire [9:0] x;  // current pixel x position: 10-bit value: 0-1023
    wire [8:0] y;  // current pixel y position:  9-bit value: 0-511
    wire animate;  // high when we're ready to animate at end of drawing
    wire collide; // collision flag
    
    //reg sq_a, sq_b, sq_c, sq_d, sq_e, sq_f, sq_g, sq_h; // registers to assign objects
    reg sq_a, sq_b, sq_c,sq_d,sq_e,sq_f; // register for rocket
    wire [11:0] sq_a_x1, sq_a_x2, sq_a_y1, sq_a_y2; // positions bits for ball
    wire [11:0] sq_b_x1, sq_b_x2, sq_b_y1, sq_b_y2; // position bits for rocket
    wire [11:0] sq_c_x1, sq_c_x2, sq_c_y1, sq_c_y2; // positions bits for decoy
    wire [11:0] sq_d_x1, sq_d_x2, sq_d_y1, sq_d_y2; // positions bits for decoy
    wire [11:0] sq_e_x1, sq_e_x2, sq_e_y1, sq_e_y2; // positions bits for decoy
    wire [11:0] sq_f_x1, sq_f_x2, sq_f_y1, sq_f_y2; // position bits for decoy
    
    wire active1;
    wire active; // active flag during game over sequence
    wire active2;
    wire [1:0] com; // bits to check rocket direction
    wire [1:0] com1; // bits to check rocket direction
    wire [1:0] com2; // bits to check rocket direction
    wire [7:0] keycode1;
    wire [7:0] keycode2;
    wire [2:0] wall1,wall2;
    assign keycode1 = keycode;
    assign keycode2 = keycode;
    
    wire player1, player2;
           
    always @(posedge CLK)
    begin
        {pix_stb, cnt} <= cnt + 16'h4000;  // divide by 4: (2^16)/4 = 0x4000
    end
    
    vga640x480 display (
        .i_clk(CLK),
        .i_pix_stb(pix_stb),
        .i_rst(mode == 2 ? &endgame : endgame[0]),
        .o_hs(VGA_HS), 
        .o_vs(VGA_VS), 
        .o_x(x), 
        .o_y(y),
        .o_animate(animate)
    ); // vga 640x480 driver
            
         
    rocket #(.P_WIDTH(RW), .P_HEIGHT(RH), .IX(RX), .IY(RY)) R1(
        .endgame(endgame|!mode),
        .i_clk(CLK), 
        .i_ani_stb(pix_stb),
        .i_animate(animate),
        .keycode(keycode),
        .o_x1(sq_b_x1),
        .o_x2(sq_b_x2),
        .o_y1(sq_b_y1),
        .o_y2(sq_b_y2),
        .active(active),
        .com(com)
        ); // rocket instance
        
      rocket2 #(.P_WIDTH(RW), .P_HEIGHT(RH), .IX(RX1), .IY(RY)) R2(
        .endgame(endgame | !mode),
        .i_clk(CLK), 
        .i_ani_stb(pix_stb),
        .i_animate(animate),
        .keycode(keycode1),
        .o_x1(sq_c_x1),
        .o_x2(sq_c_x2),
        .o_y1(sq_c_y1),
        .o_y2(sq_c_y2),
        .active(active1),
        .com(com1)
        ); // rocket instance
        
    square_4 #(.RY(RY), .RH(RH), .IX(IX), .IY(IY), .H_SIZE(B_SIZE)) b0 (
        .toggle(1 && switch == 1'b0),
        .com(com),
        .mode(mode),
        .start(active),
        .i_x1(sq_b_x1),
        .i_x2(sq_b_x2),
        .i_y1(sq_b_y1),
        .i_y2(sq_b_y2),
        .t_x1(sq_c_x1),
        .t_x2(sq_c_x2),
        .t_y1(sq_c_y1),
        .t_y2(sq_c_y2),
        .i_clk(CLK), 
        .i_ani_stb(pix_stb),
        .i_animate(animate),
        .o_x1(sq_a_x1),
        .o_x2(sq_a_x2),
        .o_y1(sq_a_y1),
        .o_y2(sq_a_y2),
        .endgame(endgame[0]),
        .score(score),
        .wall1(wall1),
        .wall2(wall2),
        .lives1(lives1),
        .lives2(lives2)
//        .RST(BTN_RST)
    ); // ball instance
    
    square1 #(.RY(RY), .RH(RH), .IX(IX), .IY(IY), .H_SIZE(B_SIZE),.wall_l(wall_l)) b1 (
        .toggle(1 && switch == 1'b1),
        .com(com),
        .mode(mode),
        .start(active),
        .i_x1(sq_b_x1),
        .i_x2(sq_b_x2),
        .i_y1(sq_b_y1),
        .i_y2(sq_b_y2),
        .t_x1(sq_c_x1),
        .t_x2(sq_c_x2),
        .t_y1(sq_c_y1),
        .t_y2(sq_c_y2),
        .i_clk(CLK), 
        .i_ani_stb(pix_stb),
        .i_animate(animate),
        .o_x1(sq_e_x1),
        .o_x2(sq_e_x2),
        .o_y1(sq_e_y1),
        .o_y2(sq_e_y2),
        .endgame(endgame[1]),
        .score(score),
        .wall1(wall1),
        .wall2(wall2),
        .lives1(lives1A)

    ); // ball instance
        square2 #(.RY(RY), .RH(RH), .IX(IX2), .IY(IY), .H_SIZE(B_SIZE),.wall_r(wall_r)) b2 (
        .toggle(1 && switch == 1'b1),
        .com(com),
        .mode(mode),
        .start(active),
        .i_x1(sq_c_x1),
        .i_x2(sq_c_x2),
        .i_y1(sq_c_y1),
        .i_y2(sq_c_y2),
        .t_x1(sq_b_x1),
        .t_x2(sq_b_x2),
        .t_y1(sq_b_y1),
        .t_y2(sq_b_y2),
        .i_clk(CLK), 
        .i_ani_stb(pix_stb),
        .i_animate(animate),
        .o_x1(sq_f_x1),
        .o_x2(sq_f_x2),
        .o_y1(sq_f_y1),
        .o_y2(sq_f_y2),
        .endgame(endgame[2]),
        .score(score),
        .wall1(wall1),
        .wall2(wall2),
        .lives2(lives2A)
    ); 

    
    always @ (*)
    begin
          sq_a = ((((x > sq_a_x1) & (y > sq_a_y1) & (x < sq_a_x2) & (y < sq_a_y2)))&& switch == 1'b0) ? 1 : 0; // draw ball edges
            sq_b = ((x > sq_b_x1) & (y > sq_b_y1) & (x < sq_b_x2) & (y < sq_b_y2)) ? 1 : 0; // draw rocket edges
            sq_c = ((x > sq_c_x1) & (y > sq_c_y1) & (x < sq_c_x2) & (y < sq_c_y2)) ? 1 : 0; // draw ball edges
            sq_d = ((x > 310) & (y > 0) & (x < 330) & (y < 480)) ? 1 : 0; // draw ball edges
            sq_e = (((x > sq_e_x1) & (y > sq_e_y1) & (x < sq_e_x2) & (y < sq_e_y2)) && switch == 1'b1) ? 1 : 0; // draw ball edges
            sq_f = (((x > sq_f_x1) & (y > sq_f_y1) & (x < sq_f_x2) & (y < sq_f_y2)) && switch == 1'b1) ? 1 : 0; // draw ball edges
            
    end
    
    always @(posedge pix_stb)
    begin
        // assign ball(s) and paddle colors

          VGA_R[3] <= ((sq_a | sq_b | sq_c | (sq_d && switch == 1'b1) | sq_e | sq_f ) && (mode == 2'b00));
          VGA_G[3] <= ((sq_a| sq_b | sq_c | (sq_d && switch == 1'b1) | sq_e | sq_f) && (mode == 2'b01)) ;
          VGA_B[3] <= (( sq_a| sq_b | sq_c | (sq_d && switch == 1'b1)| sq_e | sq_f ) && (mode == 2'b10)) ;
          VGA_R[2] <= (( sq_a |sq_b | sq_c| (sq_d && switch == 1'b1) | sq_e | sq_f) && (mode == 2'b00)) ; 
          VGA_G[2] <= (( sq_a | sq_b | sq_c |( sq_d && switch == 1'b1)| sq_e | sq_f) && (mode == 2'b01));
          VGA_B[2] <= (( sq_a| sq_b | sq_c | (sq_d && switch == 1'b1)| sq_e | sq_f) && (mode == 2'b10)) ;   
          VGA_R[1] <= (( sq_a|  sq_b | sq_c | (sq_d&& switch == 1'b1)| sq_e | sq_f) && (mode == 2'b00)) ;
          VGA_G[1] <= (( sq_a| sq_b | sq_c | (sq_d && switch == 1'b1)| sq_e | sq_f) && (mode == 2'b01)) ;
          VGA_B[1] <= (( sq_a| sq_b | sq_c | (sq_d&&switch == 1'b1)| sq_e | sq_f) && (mode == 2'b10)) ;      
          VGA_R[0] <= (( sq_a| sq_b | sq_c | (sq_d&&switch == 1'b1)| sq_e | sq_f) && (mode == 2'b00));   
          VGA_G[0] <= (( sq_a| sq_b | sq_c | (sq_d&&switch == 1'b1)| sq_e | sq_f) && (mode == 2'b01)) ;    
          VGA_B[0] <= (( sq_a| sq_b | sq_c | (sq_d && switch == 1'b1)| sq_e | sq_f) && (mode == 2'b10)) ;
    end
endmodule